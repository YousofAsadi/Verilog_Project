`timescale 1ns / 1ps

/****************************************************************************************************/
/*       __      __     _________      _       _      _________      _________      _________       */
/*       \$\    /$/    |$$$$$$$$$|    |$|     |$|    |$$$$$$$$$|    |$$$$$$$$$|    |$$$$$$$$$|      */
/*        \$\  /$/     |$|     |$|    |$|     |$|    |$|     |$|    |$|     |$|    |$|              */
/*         \$\/$/      |$|     |$|    |$|     |$|    |$|_______     |$|     |$|    |$|_____         */
/*          |$$|       |$|     |$|    |$|     |$|    |$$$$$$$$$|    |$|     |$|    |$$$$$$$|        */
/*          |$$|       |$|     |$|    |$|     |$|     _      |$|    |$|     |$|    |$|              */
/*          |$$|       |$|_____|$|    |$|_____|$|    |$|_____|$|    |$|     |$|    |$|              */
/*          |$$|       |$$$$$$$$$|    |$$$$$$$$$|    |$$$$$$$$$|    |$$$$$$$$$|    |$|              */
/*                                                                                                  */
/****************************************************************************************************/

module project_testbench;

	// Inputs
	reg x;
	reg CLK;
	reg Reset;

	// Outputs
	wire [7:0] out;

	// Instantiate the Unit Under Test (UUT)
	project uut (
		.x(x), 
		.CLK(CLK), 
		.Reset(Reset), 
		.out(out)
	);
	initial 
	begin 
	
		CLK = 1'b0;
		Reset = 1'b1;
		#15 Reset = 0;
	
	end
	
	always #5 CLK = ~CLK;
	
	initial 
	begin
		
			 x = 0;
		#10 x = 1; //
		#10 x = 1; // in sequence baraye tempreture hast
		#10 x = 1; //
		
		#10 x = 0;
		#10 x = 0;
		
		#10 x = 0; //
		#10 x = 1; // in sequence baraye humidity hast 
		#10 x = 0; //
		
		#10 x = 0;
		#10 x = 1;
		
		#10 x = 1; //
		#10 x = 0; // in sequence baraye wind hast 
		#10 x = 1; //
		
		#10 x = 1;
		#10 x = 0;
		
	end
      
endmodule

